/*
-------------------------------------------
Code  00h     defines a solid block
Codes 01h-04h define the Olin College logo
Codes 05h-1Fh define line graphics		
Codes 20h-7Eh define the ASCII characters
Code  7Fh     defines a hash pattern
Codes 80h-FFh user defined characters
-------------------------------------------
*/

module CHAR_GEN_ROM
(
pixel_clock,
address,
dataout
);

input				pixel_clock;
input [10:0]	address;
output [7:0] 	dataout;

wire [10:0] interaddr;
wire direction;
reg [7:0] data;

assign direction = 1'b1;
assign interaddr = (direction) ? {address[10:3], {3'd7 - address[2:0]}}: address;
assign dataout = (direction) ? {data[0], data[1], data[2], data[3], data[4], data[5], data[6], data[7]} : data;

always @(posedge pixel_clock) begin
	case(interaddr)
	
		//// Solid Block ////
		
		// 00h: solid block
		11'h000: data <= 8'hFF;
		11'h001: data <= 8'hFF;
		11'h002: data <= 8'hFF;
		11'h003: data <= 8'hFF;
		11'h004: data <= 8'hFF;
		11'h005: data <= 8'hFF;
		11'h006: data <= 8'hFF;
		11'h007: data <= 8'hFF;
		
		//// Logo ////
		
		// 01h: Olin "O" left half
		11'h008: data <= 8'h09;
		11'h009: data <= 8'h78;
		11'h00A: data <= 8'hF8;
		11'h00B: data <= 8'hFC;
		11'h00C: data <= 8'hFC;
		11'h00D: data <= 8'h7F;
		11'h00E: data <= 8'h0F;
		11'h00F: data <= 8'h00;
		// 02h: Olin "O" right half
		11'h010: data <= 8'hF8;
		11'h011: data <= 8'h7E;
		11'h012: data <= 8'h3F;
		11'h013: data <= 8'h1F;
		11'h014: data <= 8'h1F;
		11'h015: data <= 8'h0E;
		11'h016: data <= 8'h98;
		11'h017: data <= 8'h00;
		// 03h: Mini "OL"
		11'h018: data <= 8'h00;
		11'h019: data <= 8'h00;
		11'h01A: data <= 8'h74;
		11'h01B: data <= 8'h54;
		11'h01C: data <= 8'h54;
		11'h01D: data <= 8'h77;
		11'h01E: data <= 8'h00;
		11'h01F: data <= 8'h00;
		// 04h: Mini "IN"
		11'h020: data <= 8'h00;
		11'h021: data <= 8'h00;
		11'h022: data <= 8'h52;
		11'h023: data <= 8'h5A;
		11'h024: data <= 8'h56;
		11'h025: data <= 8'h52;
		11'h026: data <= 8'h00;
		11'h027: data <= 8'h00;
		
		//// Line Graphics ////
		
		// 05h: corner upper left
		11'h028: data <= 8'hFF;
		11'h029: data <= 8'h80;
		11'h02A: data <= 8'h80;
		11'h02B: data <= 8'h80;
		11'h02C: data <= 8'h80;
		11'h02D: data <= 8'h80;
		11'h02E: data <= 8'h80;
		11'h02F: data <= 8'h80;
		// 06h: corner upper right
		11'h030: data <= 8'hFF;
		11'h031: data <= 8'h01;
		11'h032: data <= 8'h01;
		11'h033: data <= 8'h01;
		11'h034: data <= 8'h01;
		11'h035: data <= 8'h01;
		11'h036: data <= 8'h01;
		11'h037: data <= 8'h01;
		// 07h: corner lower left
		11'h038: data <= 8'h80;
		11'h039: data <= 8'h80;
		11'h03A: data <= 8'h80;
		11'h03B: data <= 8'h80;
		11'h03C: data <= 8'h80;
		11'h03D: data <= 8'h80;
		11'h03E: data <= 8'h80;
		11'h03F: data <= 8'hFF;
		// 08h: corner lower right
		11'h040: data <= 8'h01;
		11'h041: data <= 8'h01;
		11'h042: data <= 8'h01;
		11'h043: data <= 8'h01;
		11'h044: data <= 8'h01;
		11'h045: data <= 8'h01;
		11'h046: data <= 8'h01;
		11'h047: data <= 8'hFF;
		// 09h: cross junction
		11'h048: data <= 8'h10;
		11'h049: data <= 8'h10;
		11'h04A: data <= 8'h10;
		11'h04B: data <= 8'hFF;
		11'h04C: data <= 8'h10;
		11'h04D: data <= 8'h10;
		11'h04E: data <= 8'h10;
		11'h04F: data <= 8'h10;
		// 0Ah: "T" junction
		11'h050: data <= 8'hFF;
		11'h051: data <= 8'h10;
		11'h052: data <= 8'h10;
		11'h053: data <= 8'h10;
		11'h054: data <= 8'h10;
		11'h055: data <= 8'h10;
		11'h056: data <= 8'h10;
		11'h057: data <= 8'h10;
		// 0Bh: "T" juntion rotated 90 clockwise
		11'h058: data <= 8'h01;
		11'h059: data <= 8'h01;
		11'h05A: data <= 8'h01;
		11'h05B: data <= 8'hFF;
		11'h05C: data <= 8'h01;
		11'h05D: data <= 8'h01;
		11'h05E: data <= 8'h01;
		11'h05F: data <= 8'h01;
		// 0Ch: "T" juntion rotated 180
		11'h060: data <= 8'h10;
		11'h061: data <= 8'h10;
		11'h062: data <= 8'h10;
		11'h063: data <= 8'h10;
		11'h064: data <= 8'h10;
		11'h065: data <= 8'h10;
		11'h066: data <= 8'h10;
		11'h067: data <= 8'hFF;
		// 0Dh: "T" junction rotated 270 clockwise
		11'h068: data <= 8'h80;
		11'h069: data <= 8'h80;
		11'h06A: data <= 8'h80;
		11'h06B: data <= 8'hFF;
		11'h06C: data <= 8'h80;
		11'h06D: data <= 8'h80;
		11'h06E: data <= 8'h80;
		11'h06F: data <= 8'h80;
		// 0Eh: arrow pointing right
		11'h070: data <= 8'h08;
		11'h071: data <= 8'h04;
		11'h072: data <= 8'h02;
		11'h073: data <= 8'hFF;
		11'h074: data <= 8'h02;
		11'h075: data <= 8'h04;
		11'h076: data <= 8'h08;
		11'h077: data <= 8'h00;
		// 0Fh: arrow pointing left
		11'h078: data <= 8'h10;
		11'h079: data <= 8'h20;
		11'h07A: data <= 8'h40;
		11'h07B: data <= 8'hFF;
		11'h07C: data <= 8'h40;
		11'h07D: data <= 8'h20;
		11'h07E: data <= 8'h10;
		11'h07F: data <= 8'h00;
		// 10h: first (top) horizontal line
		11'h080: data <= 8'hFF;
		11'h081: data <= 8'h00;
		11'h082: data <= 8'h00;
		11'h083: data <= 8'h00;
		11'h084: data <= 8'h00;
		11'h085: data <= 8'h00;
		11'h086: data <= 8'h00;
		11'h087: data <= 8'h00;
		// 11h: second horizontal line
		11'h088: data <= 8'h00;
		11'h089: data <= 8'hFF;
		11'h08A: data <= 8'h00;
		11'h08B: data <= 8'h00;
		11'h08C: data <= 8'h00;
		11'h08D: data <= 8'h00;
		11'h08E: data <= 8'h00;
		11'h08F: data <= 8'h00;
		// 12h: third horizontal line
		11'h090: data <= 8'h00;
		11'h091: data <= 8'h00;
		11'h092: data <= 8'hFF;
		11'h093: data <= 8'h00;
		11'h094: data <= 8'h00;
		11'h095: data <= 8'h00;
		11'h096: data <= 8'h00;
		11'h097: data <= 8'h00;
		// 13h: fourth horizontal line
		11'h098: data <= 8'h00;
		11'h099: data <= 8'h00;
		11'h09A: data <= 8'h00;
		11'h09B: data <= 8'hFF;
		11'h09C: data <= 8'h00;
		11'h09D: data <= 8'h00;
		11'h09E: data <= 8'h00;
		11'h09F: data <= 8'h00;
		// 14h: fifth horizontal line
		11'h0A0: data <= 8'h00;
		11'h0A1: data <= 8'h00;
		11'h0A2: data <= 8'h00;
		11'h0A3: data <= 8'h00;
		11'h0A4: data <= 8'hFF;
		11'h0A5: data <= 8'h00;
		11'h0A6: data <= 8'h00;
		// 15h: sixth horizontal line
		11'h0A7: data <= 8'h00;
		11'h0A8: data <= 8'h00;
		11'h0A9: data <= 8'h00;
		11'h0AA: data <= 8'h00;
		11'h0AB: data <= 8'h00;
		11'h0AC: data <= 8'h00;
		11'h0AD: data <= 8'hFF;
		11'h0AE: data <= 8'h00;
		11'h0AF: data <= 8'h00;
		// 16h: seventh horizontal line
		11'h0B0: data <= 8'h00;
		11'h0B1: data <= 8'h00;
		11'h0B2: data <= 8'h00;
		11'h0B3: data <= 8'h00;
		11'h0B4: data <= 8'h00;
		11'h0B5: data <= 8'h00;
		11'h0B6: data <= 8'hFF;
		11'h0B7: data <= 8'h00;
		// 17h: eighth (bottom) horizontal line
		11'h0B8: data <= 8'h00;
		11'h0B9: data <= 8'h00;
		11'h0BA: data <= 8'h00;
		11'h0BB: data <= 8'h00;
		11'h0BC: data <= 8'h00;
		11'h0BD: data <= 8'h00;
		11'h0BE: data <= 8'h00;
		11'h0BF: data <= 8'hFF;
		// 18h: first (left) vertical line
		11'h0C0: data <= 8'h80;
		11'h0C1: data <= 8'h80;
		11'h0C2: data <= 8'h80;
		11'h0C3: data <= 8'h80;
		11'h0C4: data <= 8'h80;
		11'h0C5: data <= 8'h80;
		11'h0C6: data <= 8'h80;
		11'h0C7: data <= 8'h80;
		// 19h: second vertical line
		11'h0C8: data <= 8'h40;
		11'h0C9: data <= 8'h40;
		11'h0CA: data <= 8'h40;
		11'h0CB: data <= 8'h40;
		11'h0CC: data <= 8'h40;
		11'h0CD: data <= 8'h40;
		11'h0CE: data <= 8'h40;
		11'h0CF: data <= 8'h40;
		// 1Ah: third vertical line
		11'h0D0: data <= 8'h20;
		11'h0D1: data <= 8'h20;
		11'h0D2: data <= 8'h20;
		11'h0D3: data <= 8'h20;
		11'h0D4: data <= 8'h20;
		11'h0D5: data <= 8'h20;
		11'h0D6: data <= 8'h20;
		11'h0D7: data <= 8'h20;
		// 1Bh: fourth vertical line
		11'h0D8: data <= 8'h10;
		11'h0D9: data <= 8'h10;
		11'h0DA: data <= 8'h10;
		11'h0DB: data <= 8'h10;
		11'h0DC: data <= 8'h10;
		11'h0DD: data <= 8'h10;
		11'h0DE: data <= 8'h10;
		11'h0DF: data <= 8'h10;
		// 1Ch: fifth vertical line
		11'h0E0: data <= 8'h08;
		11'h0E1: data <= 8'h08;
		11'h0E2: data <= 8'h08;
		11'h0E3: data <= 8'h08;
		11'h0E4: data <= 8'h08;
		11'h0E5: data <= 8'h08;
		11'h0E6: data <= 8'h08;
		11'h0E7: data <= 8'h08;
		// 1Dh: sixth vertical line
		11'h0E8: data <= 8'h04;
		11'h0E9: data <= 8'h04;
		11'h0EA: data <= 8'h04;
		11'h0EB: data <= 8'h04;
		11'h0EC: data <= 8'h04;
		11'h0ED: data <= 8'h04;
		11'h0EE: data <= 8'h04;
		11'h0EF: data <= 8'h04;
		// 1Eh: seventh vertical line
		11'h0F0: data <= 8'h02;
		11'h0F1: data <= 8'h02;
		11'h0F2: data <= 8'h02;
		11'h0F3: data <= 8'h02;
		11'h0F4: data <= 8'h02;
		11'h0F5: data <= 8'h02;
		11'h0F6: data <= 8'h02;
		11'h0F7: data <= 8'h02;
		// 1Fh: eighth (right) vertical line
		11'h0F8: data <= 8'h01;
		11'h0F9: data <= 8'h01;
		11'h0FA: data <= 8'h01;
		11'h0FB: data <= 8'h01;
		11'h0FC: data <= 8'h01;
		11'h0FD: data <= 8'h01;
		11'h0FE: data <= 8'h01;
		11'h0FF: data <= 8'h01;
		
		//// ASCII Characters ////
		
		// 20h: space
		11'h100: data <= 8'h00;
		11'h101: data <= 8'h00;
		11'h102: data <= 8'h00;
		11'h103: data <= 8'h00;
		11'h104: data <= 8'h00;
		11'h105: data <= 8'h00;
		11'h106: data <= 8'h00;
		11'h107: data <= 8'h00;
		// 21h: !
		11'h108: data <= 8'h10;
		11'h109: data <= 8'h10;
		11'h10A: data <= 8'h10;
		11'h10B: data <= 8'h10;
		11'h10C: data <= 8'h00;
		11'h10D: data <= 8'h00;
		11'h10E: data <= 8'h10;
		11'h10F: data <= 8'h00;
		// 22h: "
		11'h110: data <= 8'h28;
		11'h111: data <= 8'h28;
		11'h112: data <= 8'h28;
		11'h113: data <= 8'h00;
		11'h114: data <= 8'h00;
		11'h115: data <= 8'h00;
		11'h116: data <= 8'h00;
		11'h117: data <= 8'h00;
		// 23h: #
		11'h118: data <= 8'h28;
		11'h119: data <= 8'h28;
		11'h11A: data <= 8'h7C;
		11'h11B: data <= 8'h28;
		11'h11C: data <= 8'h7C;
		11'h11D: data <= 8'h28;
		11'h11E: data <= 8'h28;
		11'h11F: data <= 8'h00;
		// 24h: $
		11'h120: data <= 8'h10;
		11'h121: data <= 8'h3C;
		11'h122: data <= 8'h50;
		11'h123: data <= 8'h38;
		11'h124: data <= 8'h14;
		11'h125: data <= 8'h78;
		11'h126: data <= 8'h10;
		11'h127: data <= 8'h00;
		// 25h: %
		11'h128: data <= 8'h60;
		11'h129: data <= 8'h64;
		11'h12A: data <= 8'h08;
		11'h12B: data <= 8'h10;
		11'h12C: data <= 8'h20;
		11'h12D: data <= 8'h46;
		11'h12E: data <= 8'h06;
		11'h12F: data <= 8'h00;
		// 26h: &
		11'h130: data <= 8'h30;
		11'h131: data <= 8'h48;
		11'h132: data <= 8'h50;
		11'h133: data <= 8'h20;
		11'h134: data <= 8'h54;
		11'h135: data <= 8'h48;
		11'h136: data <= 8'h34;
		11'h137: data <= 8'h00;
		// 27h: '
		11'h138: data <= 8'h30;
		11'h139: data <= 8'h10;
		11'h13A: data <= 8'h20;
		11'h13B: data <= 8'h00;
		11'h13C: data <= 8'h00;
		11'h13D: data <= 8'h00;
		11'h13E: data <= 8'h00;
		11'h13F: data <= 8'h00;
		// 28h: (
		11'h140: data <= 8'h08;
		11'h141: data <= 8'h10;
		11'h142: data <= 8'h20;
		11'h143: data <= 8'h20;
		11'h144: data <= 8'h20;
		11'h145: data <= 8'h10;
		11'h146: data <= 8'h08;
		11'h147: data <= 8'h00;
		// 29h: )
		11'h148: data <= 8'h20;
		11'h149: data <= 8'h10;
		11'h14A: data <= 8'h08;
		11'h14B: data <= 8'h08;
		11'h14C: data <= 8'h08;
		11'h14D: data <= 8'h10;
		11'h14E: data <= 8'h20;
		11'h14F: data <= 8'h00;
		// 2Ah: *
		11'h150: data <= 8'h00;
		11'h151: data <= 8'h10;
		11'h152: data <= 8'h54;
		11'h153: data <= 8'h38;
		11'h154: data <= 8'h54;
		11'h155: data <= 8'h10;
		11'h156: data <= 8'h00;
		11'h157: data <= 8'h00;
		// 2Bh: +
		11'h158: data <= 8'h00;
		11'h159: data <= 8'h10;
		11'h15A: data <= 8'h10;
		11'h15B: data <= 8'h7C;
		11'h15C: data <= 8'h10;
		11'h15D: data <= 8'h10;
		11'h15E: data <= 8'h00;
		11'h15F: data <= 8'h00;
		// 2Ch: ,
		11'h160: data <= 8'h00;
		11'h161: data <= 8'h00;
		11'h162: data <= 8'h00;
		11'h163: data <= 8'h00;
		11'h164: data <= 8'h00;
		11'h165: data <= 8'h30;
		11'h166: data <= 8'h10;
		11'h167: data <= 8'h20;
		// 2Dh: -
		11'h168: data <= 8'h00;
		11'h169: data <= 8'h00;
		11'h16A: data <= 8'h00;
		11'h16B: data <= 8'h7C;
		11'h16C: data <= 8'h00;
		11'h16D: data <= 8'h00;
		11'h16E: data <= 8'h00;
		11'h16F: data <= 8'h00;
		// 2Eh: .
		11'h170: data <= 8'h00;
		11'h171: data <= 8'h00;
		11'h172: data <= 8'h00;
		11'h173: data <= 8'h00;
		11'h174: data <= 8'h00;
		11'h175: data <= 8'h30;
		11'h176: data <= 8'h30;
		11'h177: data <= 8'h00;
		// 2Fh: /
		11'h178: data <= 8'h00;
		11'h179: data <= 8'h04;
		11'h17A: data <= 8'h08;
		11'h17B: data <= 8'h10;
		11'h17C: data <= 8'h20;
		11'h17D: data <= 8'h40;
		11'h17E: data <= 8'h00;
		11'h17F: data <= 8'h00;
		// 30h: 0
		11'h180: data <= 8'h38;
		11'h181: data <= 8'h44;
		11'h182: data <= 8'h4C;
		11'h183: data <= 8'h54;
		11'h184: data <= 8'h64;
		11'h185: data <= 8'h44;
		11'h186: data <= 8'h38;
		11'h187: data <= 8'h00;
		// 31h: 1
		11'h188: data <= 8'h10;
		11'h189: data <= 8'h30;
		11'h18A: data <= 8'h10;
		11'h18B: data <= 8'h10;
		11'h18C: data <= 8'h10;
		11'h18D: data <= 8'h10;
		11'h18E: data <= 8'h38;
		11'h18F: data <= 8'h00;
		// 32h: 2
		11'h190: data <= 8'h38;
		11'h191: data <= 8'h44;
		11'h192: data <= 8'h04;
		11'h193: data <= 8'h08;
		11'h194: data <= 8'h10;
		11'h195: data <= 8'h20;
		11'h196: data <= 8'h7C;
		11'h197: data <= 8'h00;
		// 33h: 3
		11'h198: data <= 8'h7C;
		11'h199: data <= 8'h08;
		11'h19A: data <= 8'h10;
		11'h19B: data <= 8'h08;
		11'h19C: data <= 8'h04;
		11'h19D: data <= 8'h44;
		11'h19E: data <= 8'h38;
		11'h19F: data <= 8'h00;
		// 34h: 4
		11'h1A0: data <= 8'h08;
		11'h1A1: data <= 8'h18;
		11'h1A2: data <= 8'h28;
		11'h1A3: data <= 8'h48;
		11'h1A4: data <= 8'h7C;
		11'h1A5: data <= 8'h08;
		11'h1A6: data <= 8'h08;
		11'h1A7: data <= 8'h00;
		// 35h: 5
		11'h1A8: data <= 8'h7C;
		11'h1A9: data <= 8'h40;
		11'h1AA: data <= 8'h78;
		11'h1AB: data <= 8'h04;
		11'h1AC: data <= 8'h04;
		11'h1AD: data <= 8'h44;
		11'h1AE: data <= 8'h38;
		11'h1AF: data <= 8'h00;
		// 36h: 6
		11'h1B0: data <= 8'h18;
		11'h1B1: data <= 8'h20;
		11'h1B2: data <= 8'h40;
		11'h1B3: data <= 8'h78;
		11'h1B4: data <= 8'h44;
		11'h1B5: data <= 8'h44;
		11'h1B6: data <= 8'h38;
		11'h1B7: data <= 8'h00;
		// 37h: 7
		11'h1B8: data <= 8'h7C;
		11'h1B9: data <= 8'h04;
		11'h1BA: data <= 8'h08;
		11'h1BB: data <= 8'h10;
		11'h1BC: data <= 8'h20;
		11'h1BD: data <= 8'h20;
		11'h1BE: data <= 8'h20;
		11'h1BF: data <= 8'h00;
		// 38h: 8
		11'h1C0: data <= 8'h38;
		11'h1C1: data <= 8'h44;
		11'h1C2: data <= 8'h44;
		11'h1C3: data <= 8'h38;
		11'h1C4: data <= 8'h44;
		11'h1C5: data <= 8'h44;
		11'h1C6: data <= 8'h38;
		11'h1C7: data <= 8'h00;
		// 39h: 9
		11'h1C8: data <= 8'h38;
		11'h1C9: data <= 8'h44;
		11'h1CA: data <= 8'h44;
		11'h1CB: data <= 8'h3C;
		11'h1CC: data <= 8'h04;
		11'h1CD: data <= 8'h08;
		11'h1CE: data <= 8'h30;
		11'h1CF: data <= 8'h00;
		// 3Ah: :
		11'h1D0: data <= 8'h00;
		11'h1D1: data <= 8'h30;
		11'h1D2: data <= 8'h30;
		11'h1D3: data <= 8'h00;
		11'h1D4: data <= 8'h00;
		11'h1D5: data <= 8'h30;
		11'h1D6: data <= 8'h30;
		11'h1D7: data <= 8'h00;
		// 3Bh: ;
		11'h1D8: data <= 8'h00;
		11'h1D9: data <= 8'h30;
		11'h1DA: data <= 8'h30;
		11'h1DB: data <= 8'h00;
		11'h1DC: data <= 8'h00;
		11'h1DD: data <= 8'h30;
		11'h1DE: data <= 8'h10;
		11'h1DF: data <= 8'h20;
		// 3Ch: <
		11'h1E0: data <= 8'h08;
		11'h1E1: data <= 8'h10;
		11'h1E2: data <= 8'h20;
		11'h1E3: data <= 8'h40;
		11'h1E4: data <= 8'h20;
		11'h1E5: data <= 8'h10;
		11'h1E6: data <= 8'h08;
		11'h1E7: data <= 8'h00;
		// 3Dh: =
		11'h1E8: data <= 8'h00;
		11'h1E9: data <= 8'h00;
		11'h1EA: data <= 8'h7C;
		11'h1EB: data <= 8'h00;
		11'h1EC: data <= 8'h7C;
		11'h1ED: data <= 8'h00;
		11'h1EE: data <= 8'h00;
		11'h1EF: data <= 8'h00;
		// 3Eh: >
		11'h1F0: data <= 8'h20;
		11'h1F1: data <= 8'h10;
		11'h1F2: data <= 8'h08;
		11'h1F3: data <= 8'h04;
		11'h1F4: data <= 8'h08;
		11'h1F5: data <= 8'h10;
		11'h1F6: data <= 8'h20;
		11'h1F7: data <= 8'h00;
		// 3Fh: ?
		11'h1F8: data <= 8'h38;
		11'h1F9: data <= 8'h44;
		11'h1FA: data <= 8'h04;
		11'h1FB: data <= 8'h08;
		11'h1FC: data <= 8'h10;
		11'h1FD: data <= 8'h00;
		11'h1FE: data <= 8'h10;
		11'h1FF: data <= 8'h00;
		// 40h: @
		11'h200: data <= 8'h38;
		11'h201: data <= 8'h44;
		11'h202: data <= 8'h04;
		11'h203: data <= 8'h34;
		11'h204: data <= 8'h54;
		11'h205: data <= 8'h54;
		11'h206: data <= 8'h38;
		11'h207: data <= 8'h00;
		// 41h: A
		11'h208: data <= 8'h38;
		11'h209: data <= 8'h44;
		11'h20A: data <= 8'h44;
		11'h20B: data <= 8'h44;
		11'h20C: data <= 8'h7C;
		11'h20D: data <= 8'h44;
		11'h20E: data <= 8'h44;
		11'h20F: data <= 8'h00;
		// 42h: B
		11'h210: data <= 8'h78;
		11'h211: data <= 8'h44;
		11'h212: data <= 8'h44;
		11'h213: data <= 8'h78;
		11'h214: data <= 8'h44;
		11'h215: data <= 8'h44;
		11'h216: data <= 8'h78;
		11'h217: data <= 8'h00;
		// 43h: C
		11'h218: data <= 8'h38;
		11'h219: data <= 8'h44;
		11'h21A: data <= 8'h40;
		11'h21B: data <= 8'h40;
		11'h21C: data <= 8'h40;
		11'h21D: data <= 8'h44;
		11'h21E: data <= 8'h38;
		11'h21F: data <= 8'h00;
		// 44h: D
		11'h220: data <= 8'h70;
		11'h221: data <= 8'h48;
		11'h222: data <= 8'h44;
		11'h223: data <= 8'h44;
		11'h224: data <= 8'h44;
		11'h225: data <= 8'h48;
		11'h226: data <= 8'h70;
		11'h227: data <= 8'h00;
		// 45h: E
		11'h228: data <= 8'h7C;
		11'h229: data <= 8'h40;
		11'h22A: data <= 8'h40;
		11'h22B: data <= 8'h78;
		11'h22C: data <= 8'h40;
		11'h22D: data <= 8'h40;
		11'h22E: data <= 8'h7C;
		11'h22F: data <= 8'h00;
		// 46h: F
		11'h230: data <= 8'h7C;
		11'h231: data <= 8'h40;
		11'h232: data <= 8'h40;
		11'h233: data <= 8'h78;
		11'h234: data <= 8'h40;
		11'h235: data <= 8'h40;
		11'h236: data <= 8'h40;
		11'h237: data <= 8'h00;
		// 47h: G
		11'h238: data <= 8'h38;
		11'h239: data <= 8'h44;
		11'h23A: data <= 8'h40;
		11'h23B: data <= 8'h5C;
		11'h23C: data <= 8'h44;
		11'h23D: data <= 8'h44;
		11'h23E: data <= 8'h3C;
		11'h23F: data <= 8'h00;
		// 48h: H
		11'h240: data <= 8'h44;
		11'h241: data <= 8'h44;
		11'h242: data <= 8'h44;
		11'h243: data <= 8'h7C;
		11'h244: data <= 8'h44;
		11'h245: data <= 8'h44;
		11'h246: data <= 8'h44;
		11'h247: data <= 8'h00;
		// 49h: I
		11'h248: data <= 8'h38;
		11'h249: data <= 8'h10;
		11'h24A: data <= 8'h10;
		11'h24B: data <= 8'h10;
		11'h24C: data <= 8'h10;
		11'h24D: data <= 8'h10;
		11'h24E: data <= 8'h38;
		11'h24F: data <= 8'h00;
		// 4Ah: J
		11'h250: data <= 8'h1C;
		11'h251: data <= 8'h08;
		11'h252: data <= 8'h08;
		11'h253: data <= 8'h08;
		11'h254: data <= 8'h08;
		11'h255: data <= 8'h48;
		11'h256: data <= 8'h30;
		11'h257: data <= 8'h00;
		// 4Bh: K
		11'h258: data <= 8'h44;
		11'h259: data <= 8'h48;
		11'h25A: data <= 8'h50;
		11'h25B: data <= 8'h60;
		11'h25C: data <= 8'h50;
		11'h25D: data <= 8'h48;
		11'h25E: data <= 8'h44;
		11'h25F: data <= 8'h00;
		// 4Ch: L
		11'h260: data <= 8'h40;
		11'h261: data <= 8'h40;
		11'h262: data <= 8'h40;
		11'h263: data <= 8'h40;
		11'h264: data <= 8'h40;
		11'h265: data <= 8'h40;
		11'h266: data <= 8'h7C;
		11'h267: data <= 8'h00;
		// 4Dh: M
		11'h268: data <= 8'h44;
		11'h269: data <= 8'h6C;
		11'h26A: data <= 8'h54;
		11'h26B: data <= 8'h54;
		11'h26C: data <= 8'h44;
		11'h26D: data <= 8'h44;
		11'h26E: data <= 8'h44;
		11'h26F: data <= 8'h00;
		// 4Eh: N
		11'h270: data <= 8'h44;
		11'h271: data <= 8'h44;
		11'h272: data <= 8'h64;
		11'h273: data <= 8'h54;
		11'h274: data <= 8'h4C;
		11'h275: data <= 8'h44;
		11'h276: data <= 8'h44;
		11'h277: data <= 8'h00;
		// 4Fh: O
		11'h278: data <= 8'h38;
		11'h279: data <= 8'h44;
		11'h27A: data <= 8'h44;
		11'h27B: data <= 8'h44;
		11'h27C: data <= 8'h44;
		11'h27D: data <= 8'h44;
		11'h27E: data <= 8'h38;
		11'h27F: data <= 8'h00;
		// 50h: P
		11'h280: data <= 8'h78;
		11'h281: data <= 8'h44;
		11'h282: data <= 8'h44;
		11'h283: data <= 8'h78;
		11'h284: data <= 8'h40;
		11'h285: data <= 8'h40;
		11'h286: data <= 8'h40;
		11'h287: data <= 8'h00;
		// 51h: Q
		11'h288: data <= 8'h38;
		11'h289: data <= 8'h44;
		11'h28A: data <= 8'h44;
		11'h28B: data <= 8'h44;
		11'h28C: data <= 8'h54;
		11'h28D: data <= 8'h48;
		11'h28E: data <= 8'h34;
		11'h28F: data <= 8'h00;
		// 52h: R
		11'h290: data <= 8'h78;
		11'h291: data <= 8'h44;
		11'h292: data <= 8'h44;
		11'h293: data <= 8'h78;
		11'h294: data <= 8'h50;
		11'h295: data <= 8'h48;
		11'h296: data <= 8'h44;
		11'h297: data <= 8'h00;
		// 53h: S
		11'h298: data <= 8'h3C;
		11'h299: data <= 8'h40;
		11'h29A: data <= 8'h40;
		11'h29B: data <= 8'h38;
		11'h29C: data <= 8'h04;
		11'h29D: data <= 8'h04;
		11'h29E: data <= 8'h78;
		11'h29F: data <= 8'h00;
		// 54h: T
		11'h2A0: data <= 8'h7C;
		11'h2A1: data <= 8'h10;
		11'h2A2: data <= 8'h10;
		11'h2A3: data <= 8'h10;
		11'h2A4: data <= 8'h10;
		11'h2A5: data <= 8'h10;
		11'h2A6: data <= 8'h10;
		11'h2A7: data <= 8'h00;
		// 55h: U
		11'h2A8: data <= 8'h44;
		11'h2A9: data <= 8'h44;
		11'h2AA: data <= 8'h44;
		11'h2AB: data <= 8'h44;
		11'h2AC: data <= 8'h44;
		11'h2AD: data <= 8'h44;
		11'h2AE: data <= 8'h38;
		11'h2AF: data <= 8'h00;
		// 56h: V
		11'h2B0: data <= 8'h44;
		11'h2B1: data <= 8'h44;
		11'h2B2: data <= 8'h44;
		11'h2B3: data <= 8'h44;
		11'h2B4: data <= 8'h44;
		11'h2B5: data <= 8'h28;
		11'h2B6: data <= 8'h10;
		11'h2B7: data <= 8'h00;
		// 57h: W
		11'h2B8: data <= 8'h44;
		11'h2B9: data <= 8'h44;
		11'h2BA: data <= 8'h44;
		11'h2BB: data <= 8'h54;
		11'h2BC: data <= 8'h54;
		11'h2BD: data <= 8'h54;
		11'h2BE: data <= 8'h28;
		11'h2BF: data <= 8'h00;
		// 58h: X
		11'h2C0: data <= 8'h44;
		11'h2C1: data <= 8'h44;
		11'h2C2: data <= 8'h28;
		11'h2C3: data <= 8'h10;
		11'h2C4: data <= 8'h28;
		11'h2C5: data <= 8'h44;
		11'h2C6: data <= 8'h44;
		11'h2C7: data <= 8'h00;
		// 59h: Y
		11'h2C8: data <= 8'h44;
		11'h2C9: data <= 8'h44;
		11'h2CA: data <= 8'h44;
		11'h2CB: data <= 8'h28;
		11'h2CC: data <= 8'h10;
		11'h2CD: data <= 8'h10;
		11'h2CE: data <= 8'h10;
		11'h2CF: data <= 8'h00;
		// 5Ah: Z
		11'h2D0: data <= 8'h7C;
		11'h2D1: data <= 8'h04;
		11'h2D2: data <= 8'h08;
		11'h2D3: data <= 8'h10;
		11'h2D4: data <= 8'h20;
		11'h2D5: data <= 8'h40;
		11'h2D6: data <= 8'h7C;
		11'h2D7: data <= 8'h00;
		// 5Bh: [
		11'h2D8: data <= 8'h38;
		11'h2D9: data <= 8'h20;
		11'h2DA: data <= 8'h20;
		11'h2DB: data <= 8'h20;
		11'h2DC: data <= 8'h20;
		11'h2DD: data <= 8'h20;
		11'h2DE: data <= 8'h38;
		11'h2DF: data <= 8'h00;
		// 5Ch: \
		11'h2E0: data <= 8'h00;
		11'h2E1: data <= 8'h40;
		11'h2E2: data <= 8'h20;
		11'h2E3: data <= 8'h10;
		11'h2E4: data <= 8'h08;
		11'h2E5: data <= 8'h04;
		11'h2E6: data <= 8'h00;
		11'h2E7: data <= 8'h00;
		// 5Dh: ]
		11'h2E8: data <= 8'h38;
		11'h2E9: data <= 8'h08;
		11'h2EA: data <= 8'h08;
		11'h2EB: data <= 8'h08;
		11'h2EC: data <= 8'h08;
		11'h2ED: data <= 8'h08;
		11'h2EE: data <= 8'h38;
		11'h2EF: data <= 8'h00;
		// 5Eh: ^
		11'h2F0: data <= 8'h10;
		11'h2F1: data <= 8'h28;
		11'h2F2: data <= 8'h44;
		11'h2F3: data <= 8'h00;
		11'h2F4: data <= 8'h00;
		11'h2F5: data <= 8'h00;
		11'h2F6: data <= 8'h00;
		11'h2F7: data <= 8'h00;
		// 5Fh: _
		11'h2F8: data <= 8'h00;
		11'h2F9: data <= 8'h00;
		11'h2FA: data <= 8'h00;
		11'h2FB: data <= 8'h00;
		11'h2FC: data <= 8'h00;
		11'h2FD: data <= 8'h00;
		11'h2FE: data <= 8'h7C;
		11'h2FF: data <= 8'h00;
		// 60h: `
		11'h300: data <= 8'h20;
		11'h301: data <= 8'h10;
		11'h302: data <= 8'h08;
		11'h303: data <= 8'h00;
		11'h304: data <= 8'h00;
		11'h305: data <= 8'h00;
		11'h306: data <= 8'h00;
		11'h307: data <= 8'h00;
		// 61h: a
		11'h308: data <= 8'h00;
		11'h309: data <= 8'h00;
		11'h30A: data <= 8'h38;
		11'h30B: data <= 8'h04;
		11'h30C: data <= 8'h3C;
		11'h30D: data <= 8'h44;
		11'h30E: data <= 8'h3C;
		11'h30F: data <= 8'h00;
		// 62h: b
		11'h310: data <= 8'h40;
		11'h311: data <= 8'h40;
		11'h312: data <= 8'h58;
		11'h313: data <= 8'h64;
		11'h314: data <= 8'h44;
		11'h315: data <= 8'h44;
		11'h316: data <= 8'h78;
		11'h317: data <= 8'h00;
		// 63h: c
		11'h318: data <= 8'h00;
		11'h319: data <= 8'h00;
		11'h31A: data <= 8'h38;
		11'h31B: data <= 8'h40;
		11'h31C: data <= 8'h40;
		11'h31D: data <= 8'h44;
		11'h31E: data <= 8'h38;
		11'h31F: data <= 8'h00;
		// 64h: d
		11'h320: data <= 8'h04;
		11'h321: data <= 8'h04;
		11'h322: data <= 8'h34;
		11'h323: data <= 8'h4C;
		11'h324: data <= 8'h44;
		11'h325: data <= 8'h44;
		11'h326: data <= 8'h3C;
		11'h327: data <= 8'h00;
		// 65h: e
		11'h328: data <= 8'h00;
		11'h329: data <= 8'h00;
		11'h32A: data <= 8'h38;
		11'h32B: data <= 8'h44;
		11'h32C: data <= 8'h7C;
		11'h32D: data <= 8'h40;
		11'h32E: data <= 8'h38;
		11'h32F: data <= 8'h00;
		// 66h: f
		11'h330: data <= 8'h18;
		11'h331: data <= 8'h24;
		11'h332: data <= 8'h20;
		11'h333: data <= 8'h70;
		11'h334: data <= 8'h20;
		11'h335: data <= 8'h20;
		11'h336: data <= 8'h20;
		11'h337: data <= 8'h00;
		// 67h: g
		11'h338: data <= 8'h00;
		11'h339: data <= 8'h00;
		11'h33A: data <= 8'h3C;
		11'h33B: data <= 8'h44;
		11'h33C: data <= 8'h44;
		11'h33D: data <= 8'h3C;
		11'h33E: data <= 8'h04;
		11'h33F: data <= 8'h38;
		// 68h: h
		11'h340: data <= 8'h40;
		11'h341: data <= 8'h40;
		11'h342: data <= 8'h58;
		11'h343: data <= 8'h64;
		11'h344: data <= 8'h44;
		11'h345: data <= 8'h44;
		11'h346: data <= 8'h44;
		11'h347: data <= 8'h00;
		// 69h: i
		11'h348: data <= 8'h10;
		11'h349: data <= 8'h10;
		11'h34A: data <= 8'h30;
		11'h34B: data <= 8'h10;
		11'h34C: data <= 8'h10;
		11'h34D: data <= 8'h10;
		11'h34E: data <= 8'h38;
		11'h34F: data <= 8'h00;
		// 6Ah: j
		11'h350: data <= 8'h00;
		11'h351: data <= 8'h08;
		11'h352: data <= 8'h00;
		11'h353: data <= 8'h18;
		11'h354: data <= 8'h08;
		11'h355: data <= 8'h08;
		11'h356: data <= 8'h48;
		11'h357: data <= 8'h30;
		// 6Bh: k
		11'h358: data <= 8'h40;
		11'h359: data <= 8'h40;
		11'h35A: data <= 8'h48;
		11'h35B: data <= 8'h50;
		11'h35C: data <= 8'h60;
		11'h35D: data <= 8'h50;
		11'h35E: data <= 8'h48;
		11'h35F: data <= 8'h00;
		// 6Ch: l
		11'h360: data <= 8'h30;
		11'h361: data <= 8'h10;
		11'h362: data <= 8'h10;
		11'h363: data <= 8'h10;
		11'h364: data <= 8'h10;
		11'h365: data <= 8'h10;
		11'h366: data <= 8'h38;
		11'h367: data <= 8'h00;
		// 6Dh: m
		11'h368: data <= 8'h00;
		11'h369: data <= 8'h00;
		11'h36A: data <= 8'h68;
		11'h36B: data <= 8'h54;
		11'h36C: data <= 8'h54;
		11'h36D: data <= 8'h44;
		11'h36E: data <= 8'h44;
		11'h36F: data <= 8'h00;
		// 6Eh: n
		11'h370: data <= 8'h00;
		11'h371: data <= 8'h00;
		11'h372: data <= 8'h58;
		11'h373: data <= 8'h64;
		11'h374: data <= 8'h44;
		11'h375: data <= 8'h44;
		11'h376: data <= 8'h44;
		11'h377: data <= 8'h00;
		// 6Fh: o
		11'h378: data <= 8'h00;
		11'h379: data <= 8'h00;
		11'h37A: data <= 8'h38;
		11'h37B: data <= 8'h44;
		11'h37C: data <= 8'h44;
		11'h37D: data <= 8'h44;
		11'h37E: data <= 8'h38;
		11'h37F: data <= 8'h00;
		// 70h: p
		11'h380: data <= 8'h00;
		11'h381: data <= 8'h00;
		11'h382: data <= 8'h78;
		11'h383: data <= 8'h44;
		11'h384: data <= 8'h78;
		11'h385: data <= 8'h40;
		11'h386: data <= 8'h40;
		11'h387: data <= 8'h40;
		// 71h: q
		11'h388: data <= 8'h00;
		11'h389: data <= 8'h00;
		11'h38A: data <= 8'h00;
		11'h38B: data <= 8'h34;
		11'h38C: data <= 8'h4C;
		11'h38D: data <= 8'h3C;
		11'h38E: data <= 8'h04;
		11'h38F: data <= 8'h04;
		// 72h: r
		11'h390: data <= 8'h00;
		11'h391: data <= 8'h00;
		11'h392: data <= 8'h58;
		11'h393: data <= 8'h64;
		11'h394: data <= 8'h40;
		11'h395: data <= 8'h40;
		11'h396: data <= 8'h40;
		11'h397: data <= 8'h00;
		// 73h: s
		11'h398: data <= 8'h00;
		11'h399: data <= 8'h00;
		11'h39A: data <= 8'h38;
		11'h39B: data <= 8'h40;
		11'h39C: data <= 8'h38;
		11'h39D: data <= 8'h04;
		11'h39E: data <= 8'h78;
		11'h39F: data <= 8'h00;
		// 74h: t
		11'h3A0: data <= 8'h00;
		11'h3A1: data <= 8'h20;
		11'h3A2: data <= 8'h20;
		11'h3A3: data <= 8'h70;
		11'h3A4: data <= 8'h20;
		11'h3A5: data <= 8'h20;
		11'h3A6: data <= 8'h24;
		11'h3A7: data <= 8'h18;
		// 75h: u
		11'h3A8: data <= 8'h00;
		11'h3A9: data <= 8'h00;
		11'h3AA: data <= 8'h44;
		11'h3AB: data <= 8'h44;
		11'h3AC: data <= 8'h44;
		11'h3AD: data <= 8'h4C;
		11'h3AE: data <= 8'h34;
		11'h3AF: data <= 8'h00;
		// 76h: v
		11'h3B0: data <= 8'h00;
		11'h3B1: data <= 8'h00;
		11'h3B2: data <= 8'h44;
		11'h3B3: data <= 8'h44;
		11'h3B4: data <= 8'h44;
		11'h3B5: data <= 8'h28;
		11'h3B6: data <= 8'h10;
		11'h3B7: data <= 8'h00;
		// 77h: w
		11'h3B8: data <= 8'h00;
		11'h3B9: data <= 8'h00;
		11'h3BA: data <= 8'h44;
		11'h3BB: data <= 8'h44;
		11'h3BC: data <= 8'h54;
		11'h3BD: data <= 8'h54;
		11'h3BE: data <= 8'h28;
		11'h3BF: data <= 8'h00;
		// 78h: x
		11'h3C0: data <= 8'h00;
		11'h3C1: data <= 8'h00;
		11'h3C2: data <= 8'h44;
		11'h3C3: data <= 8'h28;
		11'h3C4: data <= 8'h10;
		11'h3C5: data <= 8'h28;
		11'h3C6: data <= 8'h44;
		11'h3C7: data <= 8'h00;
		// 79h: y
		11'h3C8: data <= 8'h00;
		11'h3C9: data <= 8'h00;
		11'h3CA: data <= 8'h00;
		11'h3CB: data <= 8'h44;
		11'h3CC: data <= 8'h44;
		11'h3CD: data <= 8'h3C;
		11'h3CE: data <= 8'h04;
		11'h3CF: data <= 8'h38;
		// 7Ah: z
		11'h3D0: data <= 8'h00;
		11'h3D1: data <= 8'h00;
		11'h3D2: data <= 8'h7C;
		11'h3D3: data <= 8'h08;
		11'h3D4: data <= 8'h10;
		11'h3D5: data <= 8'h20;
		11'h3D6: data <= 8'h7C;
		11'h3D7: data <= 8'h00;
		// 7Bh: {
		11'h3D8: data <= 8'h08;
		11'h3D9: data <= 8'h10;
		11'h3DA: data <= 8'h10;
		11'h3DB: data <= 8'h20;
		11'h3DC: data <= 8'h10;
		11'h3DD: data <= 8'h10;
		11'h3DE: data <= 8'h08;
		11'h3DF: data <= 8'h00;
		// 7Ch: |
		11'h3E0: data <= 8'h10;
		11'h3E1: data <= 8'h10;
		11'h3E2: data <= 8'h10;
		11'h3E3: data <= 8'h10;
		11'h3E4: data <= 8'h10;
		11'h3E5: data <= 8'h10;
		11'h3E6: data <= 8'h10;
		11'h3E7: data <= 8'h00;
		// 7Dh: }
		11'h3E8: data <= 8'h20;
		11'h3E9: data <= 8'h10;
		11'h3EA: data <= 8'h10;
		11'h3EB: data <= 8'h08;
		11'h3EC: data <= 8'h10;
		11'h3ED: data <= 8'h10;
		11'h3EE: data <= 8'h20;
		11'h3EF: data <= 8'h00;
		// 7Eh: ~
		11'h3F0: data <= 8'h00;
		11'h3F1: data <= 8'h00;
		11'h3F2: data <= 8'h60;
		11'h3F3: data <= 8'h92;
		11'h3F4: data <= 8'h0C;
		11'h3F5: data <= 8'h00;
		11'h3F6: data <= 8'h00;
		11'h3F7: data <= 8'h00;
		
		//// Hash Pattern ////
		
		// 7Fh: hash pattern
		11'h3F8: data <= 8'h55;
		11'h3F9: data <= 8'hAA;
		11'h3FA: data <= 8'h55;
		11'h3FB: data <= 8'hAA;
		11'h3FC: data <= 8'h55;
		11'h3FD: data <= 8'hAA;
		11'h3FE: data <= 8'h55;
		11'h3FF: data <= 8'hAA;
		
		//// User Defined Characters ////
		
		11'h400: data <= 8'h00;
		11'h401: data <= 8'h00;
		11'h402: data <= 8'h00;
		11'h403: data <= 8'h00;
		11'h404: data <= 8'h00;
		11'h405: data <= 8'h00;
		11'h406: data <= 8'h00;
		11'h407: data <= 8'h00;
		11'h408: data <= 8'h00;
		11'h409: data <= 8'h00;
		11'h40A: data <= 8'h00;
		11'h40B: data <= 8'h00;
		11'h40C: data <= 8'h00;
		11'h40D: data <= 8'h00;
		11'h40E: data <= 8'h00;
		11'h40F: data <= 8'h00;
		11'h410: data <= 8'h00;
		11'h411: data <= 8'h00;
		11'h412: data <= 8'h00;
		11'h413: data <= 8'h00;
		11'h414: data <= 8'h00;
		11'h415: data <= 8'h00;
		11'h416: data <= 8'h00;
		11'h417: data <= 8'h00;
		11'h418: data <= 8'h00;
		11'h419: data <= 8'h00;
		11'h41A: data <= 8'h00;
		11'h41B: data <= 8'h00;
		11'h41C: data <= 8'h00;
		11'h41D: data <= 8'h00;
		11'h41E: data <= 8'h00;
		11'h41F: data <= 8'h00;
		11'h420: data <= 8'h00;
		11'h421: data <= 8'h00;
		11'h422: data <= 8'h00;
		11'h423: data <= 8'h00;
		11'h424: data <= 8'h00;
		11'h425: data <= 8'h00;
		11'h426: data <= 8'h00;
		11'h427: data <= 8'h00;
		11'h428: data <= 8'h00;
		11'h429: data <= 8'h00;
		11'h42A: data <= 8'h00;
		11'h42B: data <= 8'h00;
		11'h42C: data <= 8'h00;
		11'h42D: data <= 8'h00;
		11'h42E: data <= 8'h00;
		11'h42F: data <= 8'h00;
		11'h430: data <= 8'h00;
		11'h431: data <= 8'h00;
		11'h432: data <= 8'h00;
		11'h433: data <= 8'h00;
		11'h434: data <= 8'h00;
		11'h435: data <= 8'h00;
		11'h436: data <= 8'h00;
		11'h437: data <= 8'h00;
		11'h438: data <= 8'h00;
		11'h439: data <= 8'h00;
		11'h43A: data <= 8'h00;
		11'h43B: data <= 8'h00;
		11'h43C: data <= 8'h00;
		11'h43D: data <= 8'h00;
		11'h43E: data <= 8'h00;
		11'h43F: data <= 8'h00;
		11'h440: data <= 8'h00;
		11'h441: data <= 8'h00;
		11'h442: data <= 8'h00;
		11'h443: data <= 8'h00;
		11'h444: data <= 8'h00;
		11'h445: data <= 8'h00;
		11'h446: data <= 8'h00;
		11'h447: data <= 8'h00;
		11'h448: data <= 8'h00;
		11'h449: data <= 8'h00;
		11'h44A: data <= 8'h00;
		11'h44B: data <= 8'h00;
		11'h44C: data <= 8'h00;
		11'h44D: data <= 8'h00;
		11'h44E: data <= 8'h00;
		11'h44F: data <= 8'h00;
		11'h450: data <= 8'h00;
		11'h451: data <= 8'h00;
		11'h452: data <= 8'h00;
		11'h453: data <= 8'h00;
		11'h454: data <= 8'h00;
		11'h455: data <= 8'h00;
		11'h456: data <= 8'h00;
		11'h457: data <= 8'h00;
		11'h458: data <= 8'h00;
		11'h459: data <= 8'h00;
		11'h45A: data <= 8'h00;
		11'h45B: data <= 8'h00;
		11'h45C: data <= 8'h00;
		11'h45D: data <= 8'h00;
		11'h45E: data <= 8'h00;
		11'h45F: data <= 8'h00;
		11'h460: data <= 8'h00;
		11'h461: data <= 8'h00;
		11'h462: data <= 8'h00;
		11'h463: data <= 8'h00;
		11'h464: data <= 8'h00;
		11'h465: data <= 8'h00;
		11'h466: data <= 8'h00;
		11'h467: data <= 8'h00;
		11'h468: data <= 8'h00;
		11'h469: data <= 8'h00;
		11'h46A: data <= 8'h00;
		11'h46B: data <= 8'h00;
		11'h46C: data <= 8'h00;
		11'h46D: data <= 8'h00;
		11'h46E: data <= 8'h00;
		11'h46F: data <= 8'h00;
		11'h470: data <= 8'h00;
		11'h471: data <= 8'h00;
		11'h472: data <= 8'h00;
		11'h473: data <= 8'h00;
		11'h474: data <= 8'h00;
		11'h475: data <= 8'h00;
		11'h476: data <= 8'h00;
		11'h477: data <= 8'h00;
		11'h478: data <= 8'h00;
		11'h479: data <= 8'h00;
		11'h47A: data <= 8'h00;
		11'h47B: data <= 8'h00;
		11'h47C: data <= 8'h00;
		11'h47D: data <= 8'h00;
		11'h47E: data <= 8'h00;
		11'h47F: data <= 8'h00;
		11'h480: data <= 8'h00;
		11'h481: data <= 8'h00;
		11'h482: data <= 8'h00;
		11'h483: data <= 8'h00;
		11'h484: data <= 8'h00;
		11'h485: data <= 8'h00;
		11'h486: data <= 8'h00;
		11'h487: data <= 8'h00;
		11'h488: data <= 8'h00;
		11'h489: data <= 8'h00;
		11'h48A: data <= 8'h00;
		11'h48B: data <= 8'h00;
		11'h48C: data <= 8'h00;
		11'h48D: data <= 8'h00;
		11'h48E: data <= 8'h00;
		11'h48F: data <= 8'h00;
		11'h490: data <= 8'h00;
		11'h491: data <= 8'h00;
		11'h492: data <= 8'h00;
		11'h493: data <= 8'h00;
		11'h494: data <= 8'h00;
		11'h495: data <= 8'h00;
		11'h496: data <= 8'h00;
		11'h497: data <= 8'h00;
		11'h498: data <= 8'h00;
		11'h499: data <= 8'h00;
		11'h49A: data <= 8'h00;
		11'h49B: data <= 8'h00;
		11'h49C: data <= 8'h00;
		11'h49D: data <= 8'h00;
		11'h49E: data <= 8'h00;
		11'h49F: data <= 8'h00;
		11'h4A0: data <= 8'h00;
		11'h4A1: data <= 8'h00;
		11'h4A2: data <= 8'h00;
		11'h4A3: data <= 8'h00;
		11'h4A4: data <= 8'h00;
		11'h4A5: data <= 8'h00;
		11'h4A6: data <= 8'h00;
		11'h4A7: data <= 8'h00;
		11'h4A8: data <= 8'h00;
		11'h4A9: data <= 8'h00;
		11'h4AA: data <= 8'h00;
		11'h4AB: data <= 8'h00;
		11'h4AC: data <= 8'h00;
		11'h4AD: data <= 8'h00;
		11'h4AE: data <= 8'h00;
		11'h4AF: data <= 8'h00;
		11'h4B0: data <= 8'h00;
		11'h4B1: data <= 8'h00;
		11'h4B2: data <= 8'h00;
		11'h4B3: data <= 8'h00;
		11'h4B4: data <= 8'h00;
		11'h4B5: data <= 8'h00;
		11'h4B6: data <= 8'h00;
		11'h4B7: data <= 8'h00;
		11'h4B8: data <= 8'h00;
		11'h4B9: data <= 8'h00;
		11'h4BA: data <= 8'h00;
		11'h4BB: data <= 8'h00;
		11'h4BC: data <= 8'h00;
		11'h4BD: data <= 8'h00;
		11'h4BE: data <= 8'h00;
		11'h4BF: data <= 8'h00;
		11'h4C0: data <= 8'h00;
		11'h4C1: data <= 8'h00;
		11'h4C2: data <= 8'h00;
		11'h4C3: data <= 8'h00;
		11'h4C4: data <= 8'h00;
		11'h4C5: data <= 8'h00;
		11'h4C6: data <= 8'h00;
		11'h4C7: data <= 8'h00;
		11'h4C8: data <= 8'h00;
		11'h4C9: data <= 8'h00;
		11'h4CA: data <= 8'h00;
		11'h4CB: data <= 8'h00;
		11'h4CC: data <= 8'h00;
		11'h4CD: data <= 8'h00;
		11'h4CE: data <= 8'h00;
		11'h4CF: data <= 8'h00;
		11'h4D0: data <= 8'h00;
		11'h4D1: data <= 8'h00;
		11'h4D2: data <= 8'h00;
		11'h4D3: data <= 8'h00;
		11'h4D4: data <= 8'h00;
		11'h4D5: data <= 8'h00;
		11'h4D6: data <= 8'h00;
		11'h4D7: data <= 8'h00;
		11'h4D8: data <= 8'h00;
		11'h4D9: data <= 8'h00;
		11'h4DA: data <= 8'h00;
		11'h4DB: data <= 8'h00;
		11'h4DC: data <= 8'h00;
		11'h4DD: data <= 8'h00;
		11'h4DE: data <= 8'h00;
		11'h4DF: data <= 8'h00;
		11'h4E0: data <= 8'h00;
		11'h4E1: data <= 8'h00;
		11'h4E2: data <= 8'h00;
		11'h4E3: data <= 8'h00;
		11'h4E4: data <= 8'h00;
		11'h4E5: data <= 8'h00;
		11'h4E6: data <= 8'h00;
		11'h4E7: data <= 8'h00;
		11'h4E8: data <= 8'h00;
		11'h4E9: data <= 8'h00;
		11'h4EA: data <= 8'h00;
		11'h4EB: data <= 8'h00;
		11'h4EC: data <= 8'h00;
		11'h4ED: data <= 8'h00;
		11'h4EE: data <= 8'h00;
		11'h4EF: data <= 8'h00;
		11'h4F0: data <= 8'h00;
		11'h4F1: data <= 8'h00;
		11'h4F2: data <= 8'h00;
		11'h4F3: data <= 8'h00;
		11'h4F4: data <= 8'h00;
		11'h4F5: data <= 8'h00;
		11'h4F6: data <= 8'h00;
		11'h4F7: data <= 8'h00;
		11'h4F8: data <= 8'h00;
		11'h4F9: data <= 8'h00;
		11'h4FA: data <= 8'h00;
		11'h4FB: data <= 8'h00;
		11'h4FC: data <= 8'h00;
		11'h4FD: data <= 8'h00;
		11'h4FE: data <= 8'h00;
		11'h4FF: data <= 8'h00;
		11'h500: data <= 8'h00;
		11'h501: data <= 8'h00;
		11'h502: data <= 8'h00;
		11'h503: data <= 8'h00;
		11'h504: data <= 8'h00;
		11'h505: data <= 8'h00;
		11'h506: data <= 8'h00;
		11'h507: data <= 8'h00;
		11'h508: data <= 8'h00;
		11'h509: data <= 8'h00;
		11'h50A: data <= 8'h00;
		11'h50B: data <= 8'h00;
		11'h50C: data <= 8'h00;
		11'h50D: data <= 8'h00;
		11'h50E: data <= 8'h00;
		11'h50F: data <= 8'h00;
		11'h510: data <= 8'h00;
		11'h511: data <= 8'h00;
		11'h512: data <= 8'h00;
		11'h513: data <= 8'h00;
		11'h514: data <= 8'h00;
		11'h515: data <= 8'h00;
		11'h516: data <= 8'h00;
		11'h517: data <= 8'h00;
		11'h518: data <= 8'h00;
		11'h519: data <= 8'h00;
		11'h51A: data <= 8'h00;
		11'h51B: data <= 8'h00;
		11'h51C: data <= 8'h00;
		11'h51D: data <= 8'h00;
		11'h51E: data <= 8'h00;
		11'h51F: data <= 8'h00;
		11'h520: data <= 8'h00;
		11'h521: data <= 8'h00;
		11'h522: data <= 8'h00;
		11'h523: data <= 8'h00;
		11'h524: data <= 8'h00;
		11'h525: data <= 8'h00;
		11'h526: data <= 8'h00;
		11'h527: data <= 8'h00;
		11'h528: data <= 8'h00;
		11'h529: data <= 8'h00;
		11'h52A: data <= 8'h00;
		11'h52B: data <= 8'h00;
		11'h52C: data <= 8'h00;
		11'h52D: data <= 8'h00;
		11'h52E: data <= 8'h00;
		11'h52F: data <= 8'h00;
		11'h530: data <= 8'h00;
		11'h531: data <= 8'h00;
		11'h532: data <= 8'h00;
		11'h533: data <= 8'h00;
		11'h534: data <= 8'h00;
		11'h535: data <= 8'h00;
		11'h536: data <= 8'h00;
		11'h537: data <= 8'h00;
		11'h538: data <= 8'h00;
		11'h539: data <= 8'h00;
		11'h53A: data <= 8'h00;
		11'h53B: data <= 8'h00;
		11'h53C: data <= 8'h00;
		11'h53D: data <= 8'h00;
		11'h53E: data <= 8'h00;
		11'h53F: data <= 8'h00;
		11'h540: data <= 8'h00;
		11'h541: data <= 8'h00;
		11'h542: data <= 8'h00;
		11'h543: data <= 8'h00;
		11'h544: data <= 8'h00;
		11'h545: data <= 8'h00;
		11'h546: data <= 8'h00;
		11'h547: data <= 8'h00;
		11'h548: data <= 8'h00;
		11'h549: data <= 8'h00;
		11'h54A: data <= 8'h00;
		11'h54B: data <= 8'h00;
		11'h54C: data <= 8'h00;
		11'h54D: data <= 8'h00;
		11'h54E: data <= 8'h00;
		11'h54F: data <= 8'h00;
		11'h550: data <= 8'h00;
		11'h551: data <= 8'h00;
		11'h552: data <= 8'h00;
		11'h553: data <= 8'h00;
		11'h554: data <= 8'h00;
		11'h555: data <= 8'h00;
		11'h556: data <= 8'h00;
		11'h557: data <= 8'h00;
		11'h558: data <= 8'h00;
		11'h559: data <= 8'h00;
		11'h55A: data <= 8'h00;
		11'h55B: data <= 8'h00;
		11'h55C: data <= 8'h00;
		11'h55D: data <= 8'h00;
		11'h55E: data <= 8'h00;
		11'h55F: data <= 8'h00;
		11'h560: data <= 8'h00;
		11'h561: data <= 8'h00;
		11'h562: data <= 8'h00;
		11'h563: data <= 8'h00;
		11'h564: data <= 8'h00;
		11'h565: data <= 8'h00;
		11'h566: data <= 8'h00;
		11'h567: data <= 8'h00;
		11'h568: data <= 8'h00;
		11'h569: data <= 8'h00;
		11'h56A: data <= 8'h00;
		11'h56B: data <= 8'h00;
		11'h56C: data <= 8'h00;
		11'h56D: data <= 8'h00;
		11'h56E: data <= 8'h00;
		11'h56F: data <= 8'h00;
		11'h570: data <= 8'h00;
		11'h571: data <= 8'h00;
		11'h572: data <= 8'h00;
		11'h573: data <= 8'h00;
		11'h574: data <= 8'h00;
		11'h575: data <= 8'h00;
		11'h576: data <= 8'h00;
		11'h577: data <= 8'h00;
		11'h578: data <= 8'h00;
		11'h579: data <= 8'h00;
		11'h57A: data <= 8'h00;
		11'h57B: data <= 8'h00;
		11'h57C: data <= 8'h00;
		11'h57D: data <= 8'h00;
		11'h57E: data <= 8'h00;
		11'h57F: data <= 8'h00;
		11'h580: data <= 8'h00;
		11'h581: data <= 8'h00;
		11'h582: data <= 8'h00;
		11'h583: data <= 8'h00;
		11'h584: data <= 8'h00;
		11'h585: data <= 8'h00;
		11'h586: data <= 8'h00;
		11'h587: data <= 8'h00;
		11'h588: data <= 8'h00;
		11'h589: data <= 8'h00;
		11'h58A: data <= 8'h00;
		11'h58B: data <= 8'h00;
		11'h58C: data <= 8'h00;
		11'h58D: data <= 8'h00;
		11'h58E: data <= 8'h00;
		11'h58F: data <= 8'h00;
		11'h590: data <= 8'h00;
		11'h591: data <= 8'h00;
		11'h592: data <= 8'h00;
		11'h593: data <= 8'h00;
		11'h594: data <= 8'h00;
		11'h595: data <= 8'h00;
		11'h596: data <= 8'h00;
		11'h597: data <= 8'h00;
		11'h598: data <= 8'h00;
		11'h599: data <= 8'h00;
		11'h59A: data <= 8'h00;
		11'h59B: data <= 8'h00;
		11'h59C: data <= 8'h00;
		11'h59D: data <= 8'h00;
		11'h59E: data <= 8'h00;
		11'h59F: data <= 8'h00;
		11'h5A0: data <= 8'h00;
		11'h5A1: data <= 8'h00;
		11'h5A2: data <= 8'h00;
		11'h5A3: data <= 8'h00;
		11'h5A4: data <= 8'h00;
		11'h5A5: data <= 8'h00;
		11'h5A6: data <= 8'h00;
		11'h5A7: data <= 8'h00;
		11'h5A8: data <= 8'h00;
		11'h5A9: data <= 8'h00;
		11'h5AA: data <= 8'h00;
		11'h5AB: data <= 8'h00;
		11'h5AC: data <= 8'h00;
		11'h5AD: data <= 8'h00;
		11'h5AE: data <= 8'h00;
		11'h5AF: data <= 8'h00;
		11'h5B0: data <= 8'h00;
		11'h5B1: data <= 8'h00;
		11'h5B2: data <= 8'h00;
		11'h5B3: data <= 8'h00;
		11'h5B4: data <= 8'h00;
		11'h5B5: data <= 8'h00;
		11'h5B6: data <= 8'h00;
		11'h5B7: data <= 8'h00;
		11'h5B8: data <= 8'h00;
		11'h5B9: data <= 8'h00;
		11'h5BA: data <= 8'h00;
		11'h5BB: data <= 8'h00;
		11'h5BC: data <= 8'h00;
		11'h5BD: data <= 8'h00;
		11'h5BE: data <= 8'h00;
		11'h5BF: data <= 8'h00;
		11'h5C0: data <= 8'h00;
		11'h5C1: data <= 8'h00;
		11'h5C2: data <= 8'h00;
		11'h5C3: data <= 8'h00;
		11'h5C4: data <= 8'h00;
		11'h5C5: data <= 8'h00;
		11'h5C6: data <= 8'h00;
		11'h5C7: data <= 8'h00;
		11'h5C8: data <= 8'h00;
		11'h5C9: data <= 8'h00;
		11'h5CA: data <= 8'h00;
		11'h5CB: data <= 8'h00;
		11'h5CC: data <= 8'h00;
		11'h5CD: data <= 8'h00;
		11'h5CE: data <= 8'h00;
		11'h5CF: data <= 8'h00;
		11'h5D0: data <= 8'h00;
		11'h5D1: data <= 8'h00;
		11'h5D2: data <= 8'h00;
		11'h5D3: data <= 8'h00;
		11'h5D4: data <= 8'h00;
		11'h5D5: data <= 8'h00;
		11'h5D6: data <= 8'h00;
		11'h5D7: data <= 8'h00;
		11'h5D8: data <= 8'h00;
		11'h5D9: data <= 8'h00;
		11'h5DA: data <= 8'h00;
		11'h5DB: data <= 8'h00;
		11'h5DC: data <= 8'h00;
		11'h5DD: data <= 8'h00;
		11'h5DE: data <= 8'h00;
		11'h5DF: data <= 8'h00;
		11'h5E0: data <= 8'h00;
		11'h5E1: data <= 8'h00;
		11'h5E2: data <= 8'h00;
		11'h5E3: data <= 8'h00;
		11'h5E4: data <= 8'h00;
		11'h5E5: data <= 8'h00;
		11'h5E6: data <= 8'h00;
		11'h5E7: data <= 8'h00;
		11'h5E8: data <= 8'h00;
		11'h5E9: data <= 8'h00;
		11'h5EA: data <= 8'h00;
		11'h5EB: data <= 8'h00;
		11'h5EC: data <= 8'h00;
		11'h5ED: data <= 8'h00;
		11'h5EE: data <= 8'h00;
		11'h5EF: data <= 8'h00;
		11'h5F0: data <= 8'h00;
		11'h5F1: data <= 8'h00;
		11'h5F2: data <= 8'h00;
		11'h5F3: data <= 8'h00;
		11'h5F4: data <= 8'h00;
		11'h5F5: data <= 8'h00;
		11'h5F6: data <= 8'h00;
		11'h5F7: data <= 8'h00;
		11'h5F8: data <= 8'h00;
		11'h5F9: data <= 8'h00;
		11'h5FA: data <= 8'h00;
		11'h5FB: data <= 8'h00;
		11'h5FC: data <= 8'h00;
		11'h5FD: data <= 8'h00;
		11'h5FE: data <= 8'h00;
		11'h5FF: data <= 8'h00;
		11'h600: data <= 8'h00;
		11'h601: data <= 8'h00;
		11'h602: data <= 8'h00;
		11'h603: data <= 8'h00;
		11'h604: data <= 8'h00;
		11'h605: data <= 8'h00;
		11'h606: data <= 8'h00;
		11'h607: data <= 8'h00;
		11'h608: data <= 8'h00;
		11'h609: data <= 8'h00;
		11'h60A: data <= 8'h00;
		11'h60B: data <= 8'h00;
		11'h60C: data <= 8'h00;
		11'h60D: data <= 8'h00;
		11'h60E: data <= 8'h00;
		11'h60F: data <= 8'h00;
		11'h610: data <= 8'h00;
		11'h611: data <= 8'h00;
		11'h612: data <= 8'h00;
		11'h613: data <= 8'h00;
		11'h614: data <= 8'h00;
		11'h615: data <= 8'h00;
		11'h616: data <= 8'h00;
		11'h617: data <= 8'h00;
		11'h618: data <= 8'h00;
		11'h619: data <= 8'h00;
		11'h61A: data <= 8'h00;
		11'h61B: data <= 8'h00;
		11'h61C: data <= 8'h00;
		11'h61D: data <= 8'h00;
		11'h61E: data <= 8'h00;
		11'h61F: data <= 8'h00;
		11'h620: data <= 8'h00;
		11'h621: data <= 8'h00;
		11'h622: data <= 8'h00;
		11'h623: data <= 8'h00;
		11'h624: data <= 8'h00;
		11'h625: data <= 8'h00;
		11'h626: data <= 8'h00;
		11'h627: data <= 8'h00;
		11'h628: data <= 8'h00;
		11'h629: data <= 8'h00;
		11'h62A: data <= 8'h00;
		11'h62B: data <= 8'h00;
		11'h62C: data <= 8'h00;
		11'h62D: data <= 8'h00;
		11'h62E: data <= 8'h00;
		11'h62F: data <= 8'h00;
		11'h630: data <= 8'h00;
		11'h631: data <= 8'h00;
		11'h632: data <= 8'h00;
		11'h633: data <= 8'h00;
		11'h634: data <= 8'h00;
		11'h635: data <= 8'h00;
		11'h636: data <= 8'h00;
		11'h637: data <= 8'h00;
		11'h638: data <= 8'h00;
		11'h639: data <= 8'h00;
		11'h63A: data <= 8'h00;
		11'h63B: data <= 8'h00;
		11'h63C: data <= 8'h00;
		11'h63D: data <= 8'h00;
		11'h63E: data <= 8'h00;
		11'h63F: data <= 8'h00;
		11'h640: data <= 8'h00;
		11'h641: data <= 8'h00;
		11'h642: data <= 8'h00;
		11'h643: data <= 8'h00;
		11'h644: data <= 8'h00;
		11'h645: data <= 8'h00;
		11'h646: data <= 8'h00;
		11'h647: data <= 8'h00;
		11'h648: data <= 8'h00;
		11'h649: data <= 8'h00;
		11'h64A: data <= 8'h00;
		11'h64B: data <= 8'h00;
		11'h64C: data <= 8'h00;
		11'h64D: data <= 8'h00;
		11'h64E: data <= 8'h00;
		11'h64F: data <= 8'h00;
		11'h650: data <= 8'h00;
		11'h651: data <= 8'h00;
		11'h652: data <= 8'h00;
		11'h653: data <= 8'h00;
		11'h654: data <= 8'h00;
		11'h655: data <= 8'h00;
		11'h656: data <= 8'h00;
		11'h657: data <= 8'h00;
		11'h658: data <= 8'h00;
		11'h659: data <= 8'h00;
		11'h65A: data <= 8'h00;
		11'h65B: data <= 8'h00;
		11'h65C: data <= 8'h00;
		11'h65D: data <= 8'h00;
		11'h65E: data <= 8'h00;
		11'h65F: data <= 8'h00;
		11'h660: data <= 8'h00;
		11'h661: data <= 8'h00;
		11'h662: data <= 8'h00;
		11'h663: data <= 8'h00;
		11'h664: data <= 8'h00;
		11'h665: data <= 8'h00;
		11'h666: data <= 8'h00;
		11'h667: data <= 8'h00;
		11'h668: data <= 8'h00;
		11'h669: data <= 8'h00;
		11'h66A: data <= 8'h00;
		11'h66B: data <= 8'h00;
		11'h66C: data <= 8'h00;
		11'h66D: data <= 8'h00;
		11'h66E: data <= 8'h00;
		11'h66F: data <= 8'h00;
		11'h670: data <= 8'h00;
		11'h671: data <= 8'h00;
		11'h672: data <= 8'h00;
		11'h673: data <= 8'h00;
		11'h674: data <= 8'h00;
		11'h675: data <= 8'h00;
		11'h676: data <= 8'h00;
		11'h677: data <= 8'h00;
		11'h678: data <= 8'h00;
		11'h679: data <= 8'h00;
		11'h67A: data <= 8'h00;
		11'h67B: data <= 8'h00;
		11'h67C: data <= 8'h00;
		11'h67D: data <= 8'h00;
		11'h67E: data <= 8'h00;
		11'h67F: data <= 8'h00;
		11'h680: data <= 8'h00;
		11'h681: data <= 8'h00;
		11'h682: data <= 8'h00;
		11'h683: data <= 8'h00;
		11'h684: data <= 8'h00;
		11'h685: data <= 8'h00;
		11'h686: data <= 8'h00;
		11'h687: data <= 8'h00;
		11'h688: data <= 8'h00;
		11'h689: data <= 8'h00;
		11'h68A: data <= 8'h00;
		11'h68B: data <= 8'h00;
		11'h68C: data <= 8'h00;
		11'h68D: data <= 8'h00;
		11'h68E: data <= 8'h00;
		11'h68F: data <= 8'h00;
		11'h690: data <= 8'h00;
		11'h691: data <= 8'h00;
		11'h692: data <= 8'h00;
		11'h693: data <= 8'h00;
		11'h694: data <= 8'h00;
		11'h695: data <= 8'h00;
		11'h696: data <= 8'h00;
		11'h697: data <= 8'h00;
		11'h698: data <= 8'h00;
		11'h699: data <= 8'h00;
		11'h69A: data <= 8'h00;
		11'h69B: data <= 8'h00;
		11'h69C: data <= 8'h00;
		11'h69D: data <= 8'h00;
		11'h69E: data <= 8'h00;
		11'h69F: data <= 8'h00;
		11'h6A0: data <= 8'h00;
		11'h6A1: data <= 8'h00;
		11'h6A2: data <= 8'h00;
		11'h6A3: data <= 8'h00;
		11'h6A4: data <= 8'h00;
		11'h6A5: data <= 8'h00;
		11'h6A6: data <= 8'h00;
		11'h6A7: data <= 8'h00;
		11'h6A8: data <= 8'h00;
		11'h6A9: data <= 8'h00;
		11'h6AA: data <= 8'h00;
		11'h6AB: data <= 8'h00;
		11'h6AC: data <= 8'h00;
		11'h6AD: data <= 8'h00;
		11'h6AE: data <= 8'h00;
		11'h6AF: data <= 8'h00;
		11'h6B0: data <= 8'h00;
		11'h6B1: data <= 8'h00;
		11'h6B2: data <= 8'h00;
		11'h6B3: data <= 8'h00;
		11'h6B4: data <= 8'h00;
		11'h6B5: data <= 8'h00;
		11'h6B6: data <= 8'h00;
		11'h6B7: data <= 8'h00;
		11'h6B8: data <= 8'h00;
		11'h6B9: data <= 8'h00;
		11'h6BA: data <= 8'h00;
		11'h6BB: data <= 8'h00;
		11'h6BC: data <= 8'h00;
		11'h6BD: data <= 8'h00;
		11'h6BE: data <= 8'h00;
		11'h6BF: data <= 8'h00;
		11'h6C0: data <= 8'h00;
		11'h6C1: data <= 8'h00;
		11'h6C2: data <= 8'h00;
		11'h6C3: data <= 8'h00;
		11'h6C4: data <= 8'h00;
		11'h6C5: data <= 8'h00;
		11'h6C6: data <= 8'h00;
		11'h6C7: data <= 8'h00;
		11'h6C8: data <= 8'h00;
		11'h6C9: data <= 8'h00;
		11'h6CA: data <= 8'h00;
		11'h6CB: data <= 8'h00;
		11'h6CC: data <= 8'h00;
		11'h6CD: data <= 8'h00;
		11'h6CE: data <= 8'h00;
		11'h6CF: data <= 8'h00;
		11'h6D0: data <= 8'h00;
		11'h6D1: data <= 8'h00;
		11'h6D2: data <= 8'h00;
		11'h6D3: data <= 8'h00;
		11'h6D4: data <= 8'h00;
		11'h6D5: data <= 8'h00;
		11'h6D6: data <= 8'h00;
		11'h6D7: data <= 8'h00;
		11'h6D8: data <= 8'h00;
		11'h6D9: data <= 8'h00;
		11'h6DA: data <= 8'h00;
		11'h6DB: data <= 8'h00;
		11'h6DC: data <= 8'h00;
		11'h6DD: data <= 8'h00;
		11'h6DE: data <= 8'h00;
		11'h6DF: data <= 8'h00;
		11'h6E0: data <= 8'h00;
		11'h6E1: data <= 8'h00;
		11'h6E2: data <= 8'h00;
		11'h6E3: data <= 8'h00;
		11'h6E4: data <= 8'h00;
		11'h6E5: data <= 8'h00;
		11'h6E6: data <= 8'h00;
		11'h6E7: data <= 8'h00;
		11'h6E8: data <= 8'h00;
		11'h6E9: data <= 8'h00;
		11'h6EA: data <= 8'h00;
		11'h6EB: data <= 8'h00;
		11'h6EC: data <= 8'h00;
		11'h6ED: data <= 8'h00;
		11'h6EE: data <= 8'h00;
		11'h6EF: data <= 8'h00;
		11'h6F0: data <= 8'h00;
		11'h6F1: data <= 8'h00;
		11'h6F2: data <= 8'h00;
		11'h6F3: data <= 8'h00;
		11'h6F4: data <= 8'h00;
		11'h6F5: data <= 8'h00;
		11'h6F6: data <= 8'h00;
		11'h6F7: data <= 8'h00;
		11'h6F8: data <= 8'h00;
		11'h6F9: data <= 8'h00;
		11'h6FA: data <= 8'h00;
		11'h6FB: data <= 8'h00;
		11'h6FC: data <= 8'h00;
		11'h6FD: data <= 8'h00;
		11'h6FE: data <= 8'h00;
		11'h6FF: data <= 8'h00;
		11'h700: data <= 8'h00;
		11'h701: data <= 8'h00;
		11'h702: data <= 8'h00;
		11'h703: data <= 8'h00;
		11'h704: data <= 8'h00;
		11'h705: data <= 8'h00;
		11'h706: data <= 8'h00;
		11'h707: data <= 8'h00;
		11'h708: data <= 8'h00;
		11'h709: data <= 8'h00;
		11'h70A: data <= 8'h00;
		11'h70B: data <= 8'h00;
		11'h70C: data <= 8'h00;
		11'h70D: data <= 8'h00;
		11'h70E: data <= 8'h00;
		11'h70F: data <= 8'h00;
		11'h710: data <= 8'h00;
		11'h711: data <= 8'h00;
		11'h712: data <= 8'h00;
		11'h713: data <= 8'h00;
		11'h714: data <= 8'h00;
		11'h715: data <= 8'h00;
		11'h716: data <= 8'h00;
		11'h717: data <= 8'h00;
		11'h718: data <= 8'h00;
		11'h719: data <= 8'h00;
		11'h71A: data <= 8'h00;
		11'h71B: data <= 8'h00;
		11'h71C: data <= 8'h00;
		11'h71D: data <= 8'h00;
		11'h71E: data <= 8'h00;
		11'h71F: data <= 8'h00;
		11'h720: data <= 8'h00;
		11'h721: data <= 8'h00;
		11'h722: data <= 8'h00;
		11'h723: data <= 8'h00;
		11'h724: data <= 8'h00;
		11'h725: data <= 8'h00;
		11'h726: data <= 8'h00;
		11'h727: data <= 8'h00;
		11'h728: data <= 8'h00;
		11'h729: data <= 8'h00;
		11'h72A: data <= 8'h00;
		11'h72B: data <= 8'h00;
		11'h72C: data <= 8'h00;
		11'h72D: data <= 8'h00;
		11'h72E: data <= 8'h00;
		11'h72F: data <= 8'h00;
		11'h730: data <= 8'h00;
		11'h731: data <= 8'h00;
		11'h732: data <= 8'h00;
		11'h733: data <= 8'h00;
		11'h734: data <= 8'h00;
		11'h735: data <= 8'h00;
		11'h736: data <= 8'h00;
		11'h737: data <= 8'h00;
		11'h738: data <= 8'h00;
		11'h739: data <= 8'h00;
		11'h73A: data <= 8'h00;
		11'h73B: data <= 8'h00;
		11'h73C: data <= 8'h00;
		11'h73D: data <= 8'h00;
		11'h73E: data <= 8'h00;
		11'h73F: data <= 8'h00;
		11'h740: data <= 8'h00;
		11'h741: data <= 8'h00;
		11'h742: data <= 8'h00;
		11'h743: data <= 8'h00;
		11'h744: data <= 8'h00;
		11'h745: data <= 8'h00;
		11'h746: data <= 8'h00;
		11'h747: data <= 8'h00;
		11'h748: data <= 8'h00;
		11'h749: data <= 8'h00;
		11'h74A: data <= 8'h00;
		11'h74B: data <= 8'h00;
		11'h74C: data <= 8'h00;
		11'h74D: data <= 8'h00;
		11'h74E: data <= 8'h00;
		11'h74F: data <= 8'h00;
		11'h750: data <= 8'h00;
		11'h751: data <= 8'h00;
		11'h752: data <= 8'h00;
		11'h753: data <= 8'h00;
		11'h754: data <= 8'h00;
		11'h755: data <= 8'h00;
		11'h756: data <= 8'h00;
		11'h757: data <= 8'h00;
		11'h758: data <= 8'h00;
		11'h759: data <= 8'h00;
		11'h75A: data <= 8'h00;
		11'h75B: data <= 8'h00;
		11'h75C: data <= 8'h00;
		11'h75D: data <= 8'h00;
		11'h75E: data <= 8'h00;
		11'h75F: data <= 8'h00;
		11'h760: data <= 8'h00;
		11'h761: data <= 8'h00;
		11'h762: data <= 8'h00;
		11'h763: data <= 8'h00;
		11'h764: data <= 8'h00;
		11'h765: data <= 8'h00;
		11'h766: data <= 8'h00;
		11'h767: data <= 8'h00;
		11'h768: data <= 8'h00;
		11'h769: data <= 8'h00;
		11'h76A: data <= 8'h00;
		11'h76B: data <= 8'h00;
		11'h76C: data <= 8'h00;
		11'h76D: data <= 8'h00;
		11'h76E: data <= 8'h00;
		11'h76F: data <= 8'h00;
		11'h770: data <= 8'h00;
		11'h771: data <= 8'h00;
		11'h772: data <= 8'h00;
		11'h773: data <= 8'h00;
		11'h774: data <= 8'h00;
		11'h775: data <= 8'h00;
		11'h776: data <= 8'h00;
		11'h777: data <= 8'h00;
		11'h778: data <= 8'h00;
		11'h779: data <= 8'h00;
		11'h77A: data <= 8'h00;
		11'h77B: data <= 8'h00;
		11'h77C: data <= 8'h00;
		11'h77D: data <= 8'h00;
		11'h77E: data <= 8'h00;
		11'h77F: data <= 8'h00;
		11'h780: data <= 8'h00;
		11'h781: data <= 8'h00;
		11'h782: data <= 8'h00;
		11'h783: data <= 8'h00;
		11'h784: data <= 8'h00;
		11'h785: data <= 8'h00;
		11'h786: data <= 8'h00;
		11'h787: data <= 8'h00;
		11'h788: data <= 8'h00;
		11'h789: data <= 8'h00;
		11'h78A: data <= 8'h00;
		11'h78B: data <= 8'h00;
		11'h78C: data <= 8'h00;
		11'h78D: data <= 8'h00;
		11'h78E: data <= 8'h00;
		11'h78F: data <= 8'h00;
		11'h790: data <= 8'h00;
		11'h791: data <= 8'h00;
		11'h792: data <= 8'h00;
		11'h793: data <= 8'h00;
		11'h794: data <= 8'h00;
		11'h795: data <= 8'h00;
		11'h796: data <= 8'h00;
		11'h797: data <= 8'h00;
		11'h798: data <= 8'h00;
		11'h799: data <= 8'h00;
		11'h79A: data <= 8'h00;
		11'h79B: data <= 8'h00;
		11'h79C: data <= 8'h00;
		11'h79D: data <= 8'h00;
		11'h79E: data <= 8'h00;
		11'h79F: data <= 8'h00;
		11'h7A0: data <= 8'h00;
		11'h7A1: data <= 8'h00;
		11'h7A2: data <= 8'h00;
		11'h7A3: data <= 8'h00;
		11'h7A4: data <= 8'h00;
		11'h7A5: data <= 8'h00;
		11'h7A6: data <= 8'h00;
		11'h7A7: data <= 8'h00;
		11'h7A8: data <= 8'h00;
		11'h7A9: data <= 8'h00;
		11'h7AA: data <= 8'h00;
		11'h7AB: data <= 8'h00;
		11'h7AC: data <= 8'h00;
		11'h7AD: data <= 8'h00;
		11'h7AE: data <= 8'h00;
		11'h7AF: data <= 8'h00;
		11'h7B0: data <= 8'h00;
		11'h7B1: data <= 8'h00;
		11'h7B2: data <= 8'h00;
		11'h7B3: data <= 8'h00;
		11'h7B4: data <= 8'h00;
		11'h7B5: data <= 8'h00;
		11'h7B6: data <= 8'h00;
		11'h7B7: data <= 8'h00;
		11'h7B8: data <= 8'h00;
		11'h7B9: data <= 8'h00;
		11'h7BA: data <= 8'h00;
		11'h7BB: data <= 8'h00;
		11'h7BC: data <= 8'h00;
		11'h7BD: data <= 8'h00;
		11'h7BE: data <= 8'h00;
		11'h7BF: data <= 8'h00;
		11'h7C0: data <= 8'h00;
		11'h7C1: data <= 8'h00;
		11'h7C2: data <= 8'h00;
		11'h7C3: data <= 8'h00;
		11'h7C4: data <= 8'h00;
		11'h7C5: data <= 8'h00;
		11'h7C6: data <= 8'h00;
		11'h7C7: data <= 8'h00;
		11'h7C8: data <= 8'h00;
		11'h7C9: data <= 8'h00;
		11'h7CA: data <= 8'h00;
		11'h7CB: data <= 8'h00;
		11'h7CC: data <= 8'h00;
		11'h7CD: data <= 8'h00;
		11'h7CE: data <= 8'h00;
		11'h7CF: data <= 8'h00;
		11'h7D0: data <= 8'h00;
		11'h7D1: data <= 8'h00;
		11'h7D2: data <= 8'h00;
		11'h7D3: data <= 8'h00;
		11'h7D4: data <= 8'h00;
		11'h7D5: data <= 8'h00;
		11'h7D6: data <= 8'h00;
		11'h7D7: data <= 8'h00;
		11'h7D8: data <= 8'h00;
		11'h7D9: data <= 8'h00;
		11'h7DA: data <= 8'h00;
		11'h7DB: data <= 8'h00;
		11'h7DC: data <= 8'h00;
		11'h7DD: data <= 8'h00;
		11'h7DE: data <= 8'h00;
		11'h7DF: data <= 8'h00;
		11'h7E0: data <= 8'h00;
		11'h7E1: data <= 8'h00;
		11'h7E2: data <= 8'h00;
		11'h7E3: data <= 8'h00;
		11'h7E4: data <= 8'h00;
		11'h7E5: data <= 8'h00;
		11'h7E6: data <= 8'h00;
		11'h7E7: data <= 8'h00;
		11'h7E8: data <= 8'h00;
		11'h7E9: data <= 8'h00;
		11'h7EA: data <= 8'h00;
		11'h7EB: data <= 8'h00;
		11'h7EC: data <= 8'h00;
		11'h7ED: data <= 8'h00;
		11'h7EE: data <= 8'h00;
		11'h7EF: data <= 8'h00;
		11'h7F0: data <= 8'h00;
		11'h7F1: data <= 8'h00;
		11'h7F2: data <= 8'h00;
		11'h7F3: data <= 8'h00;
		11'h7F4: data <= 8'h00;
		11'h7F5: data <= 8'h00;
		11'h7F6: data <= 8'h00;
		11'h7F7: data <= 8'h00;
		11'h7F8: data <= 8'h00;
		11'h7F9: data <= 8'h00;
		11'h7FA: data <= 8'h00;
		11'h7FB: data <= 8'h00;
		11'h7FC: data <= 8'h00;
		11'h7FD: data <= 8'h00;
		11'h7FE: data <= 8'h00;
		11'h7FF: data <= 8'h00;
	endcase                              
end

endmodule //CHAR_GEN_ROM




